-- top level entity
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity astrocam is
  port (
    clk : in std_logic;
    rst : in std_logic
  );
end astrocam;

architecture structural of astrocam is

begin

end architecture;